module webview

#flag windows -L@VMODROOT/webview/webview2/build/native/x64 -lWebView2Loader.dll
#flag windows -lole32 -lshell32 -lshlwapi -luser32
#flag windows -I @VMODROOT/webview/webview2/build/native/include
#flag -static

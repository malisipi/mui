module webview

#pkgconfig gtk+-3.0
#pkgconfig webkit2gtk-4.0

module mui

pub fn C.emscripten_run_script(a &char)
pub fn C.emscripten_run_script_string(a &char) &char
//pub fn C.emscripten_run_async_script(a &char)

const (
    text_cursor="|"
    os_font="noto.ttf"
)

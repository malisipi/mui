module window

fn C.gtk_widget_hide(win voidptr)
fn C.gtk_widget_show(win voidptr)
fn C.putenv(&char) int

module mui

import os

const(
	narrator_vbs=os.temp_dir()+"/mui_speak.vbs"
)

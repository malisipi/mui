module mui

pub fn C.emscripten_run_script(&char)
pub fn C.emscripten_run_script_string(&char) &char
pub fn C.emscripten_sleep(int)
//pub fn C.emscripten_run_async_script(&char)

const (
    text_cursor="|"
    os_font="noto.ttf"
)

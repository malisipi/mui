module mui

import os.font

const text_cursor="|"
const os_font=font.default()

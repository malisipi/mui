module mui

fn C.mui_get_regedit_dword(&u16, &u16) &u16
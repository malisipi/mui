module window

fn C.FreeConsole()
fn C.AllocConsole()
fn C.GetConsoleWindow() voidptr
fn C.ShowWindow(voidptr, bool)

module mui

const (
    text_cursor="│"
)

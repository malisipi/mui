module mui

import os.font

const (
    text_cursor="|"
    os_font=font.default()
)

module mui

const (
	hiragana_list={
		"んあ":"な", //fix na/ni/nu/ne/no letters
		"んい":"に",
		"んう":"ぬ",
		"んえ":"ね",
		"んお":"の",

		"a":"あ",
		"i":"い",
		"u":"う",
		"e":"え",
		"o":"お",
		"n":"ん",
		"ya":"ゃ",
		"yu":"ゅ",
		"yo":"ょ",
		"va":"ゎ",
		"ka":"か",
		"ki":"き",
		"ku":"く",
		"ke":"け",
		"ko":"こ",
		"sa":"さ",
		"su":"す",
		"se":"せ",
		"so":"そ",
		"ta":"た",
		"chi":"ち",
		"tsu":"つ",
		"te":"て",
		"to":"と",
		"na":"な",
		"ni":"に",
		"nu":"ぬ",
		"ne":"ね",
		"no":"の",
		"ha":"は",
		"hi":"ひ",
		"fu":"ふ",
		"he":"へ",
		"ho":"ほ",
		"ma":"ま",
		"mi":"み",
		"mu":"む",
		"me":"め",
		"mo":"も",
		"ra":"ら",
		"ri":"り",
		"ru":"る",
		"re":"れ",
		"ro":"ろ",
		"vi":"ゐ",
		"ve":"ゑ",
		"vo":"を",
		"ga":"が",
		"gi":"ぎ",
		"gu":"ぐ",
		"ge":"げ",
		"go":"ご",
		"za":"ざ",
		"ji":"じ",
		"zu":"ず",
		"ze":"ぜ",
		"zo":"ぞ",
		"da":"だ",
		"ci":"ぢ",
		"de":"で",
		"do":"ど",
		"ca":"ぢゃ",
		"cu":"ぢゅ",
		"co":"ぢょ",
		"ba":"ば",
		"bi":"び",
		"bu":"ぶ",
		"be":"べ",
		"bo":"ぼ",
		"pa":"ぱ",
		"pi":"ぴ",
		"pu":"ぷ",
		"pe":"ぺ",
		"po":"ぽ",
		"dzu":"づ",
		"shi":"し",
		"kya":"きゃ",
		"kyu":"きゅ",
		"kyo":"きょ",
		"kva":"くゎ",
		"sha":"しゃ",
		"shu":"しゅ",
		"sho":"しょ",
		"cha":"ちゃ",
		"chu":"ちゅ",
		"cho":"ちょ",
		"nya":"にゃ",
		"nyu":"にゅ",
		"nyo":"にょ",
		"hya":"ひゃ",
		"hyu":"ひゅ",
		"hyo":"ひょ",
		"mya":"みゃ",
		"myu":"みゅ",
		"myo":"みょ",
		"rya":"りゃ",
		"ryu":"りゅ",
		"ryo":"りょ",
		"gya":"ぎゃ",
		"gyu":"ぎゅ",
		"gyo":"ぎょ",
		"gva":"ぐゎ",
		"bya":"びゃ",
		"byu":"びゅ",
		"byo":"びょ",
		"pya":"ぴゃ",
		"pyu":"ぴゅ",
		"pyo":"ぴょ"
	}
	hiragana_keys=unsafe { hiragana_list.keys().clone().reverse() }
)

fn replace_romanji_with_hiragana (romanji string) string {
	mut hiragana := romanji.clone()
	for hkey in hiragana_keys {
		hiragana = hiragana.replace(hkey, hiragana_list[hkey])
	}
	return hiragana
}
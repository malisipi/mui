module mui

fn C.GetKeyState(key int) bool
module mui

fn about_dialog(event_details EventDetails, mut app &Window, app_data voidptr){
	messagebox("MUI","MUI -  1.0.0\n* TinyFileDialogs: 3.8.8","ok","info")
}
